module CharGenSlave(dat_i, dat_o, ack_o, adr_i, cyc_i,
    err_o, rty_o, sel_i, stb_i, we_i,
    clk_bus, rst_bus, hdata, vdata, dvi_red, dvi_blue, dvi_green,
    de_hp, de_vp, de_svp, de_valid, de_ascii);

input wire clk_bus;
input wire rst_bus;

// ----------- system bus slave interface ---------


input wire [31:0] dat_i;
output wire [31:0] dat_o;
output wire ack_o;
input wire [31:0] adr_i;
input wire cyc_i;
output wire err_o;
output wire rty_o;
input wire [3:0] sel_i;
input wire stb_i;
input wire we_i;

// ----------------- video io ------------

input wire [11:0] hdata;
input wire [11:0] vdata;


output wire [2:0] dvi_red;
output wire [2:0] dvi_green;
output wire [1:0] dvi_blue;

// for debugging
output wire [6:0] de_hp;
output wire [6:0] de_vp;
output wire [6:0] de_svp;
output wire de_valid;
output wire [7:0] de_ascii;

reg [31:0] stored_dat;
reg [6:0] svp; // the first row number
reg [6:0] hp;
reg [6:0] vp;
wire [6:0] next_svp;
wire [6:0] next_hp;
wire [6:0] next_vp;
wire next_full;

reg full;
integer i;
integer j;

wire [6:0] char_hdata;
wire [6:0] char_vdata;
wire [2:0] char_ih;
wire [2:0] char_iv;
wire [7:0] char_code;
wire pixel;
wire valid; // the position has been occupied by a character
wire painted; // the position has pixel

reg [7:0] char_ram[74:0][99:0];
wire [7:0] next_char_ram[74:0][99:0];
// reg [63:0] font_rom[0:127];
parameter [128 * 64 - 1 : 0] font_rom = {
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00111011,8'b01101110,
    8'b00000000,8'b00000111,8'b00001100,8'b00001100,8'b00111000,8'b00001100,8'b00001100,8'b00000111,
    8'b00000000,8'b00011000,8'b00011000,8'b00011000,8'b00000000,8'b00011000,8'b00011000,8'b00011000,
    8'b00000000,8'b00111000,8'b00001100,8'b00001100,8'b00000111,8'b00001100,8'b00001100,8'b00111000,
    8'b00000000,8'b00111111,8'b00100110,8'b00001100,8'b00011001,8'b00111111,8'b00000000,8'b00000000,
    8'b00011111,8'b00110000,8'b00111110,8'b00110011,8'b00110011,8'b00110011,8'b00000000,8'b00000000,
    8'b00000000,8'b01100011,8'b00110110,8'b00011100,8'b00110110,8'b01100011,8'b00000000,8'b00000000,
    8'b00000000,8'b00110110,8'b01111111,8'b01111111,8'b01101011,8'b01100011,8'b00000000,8'b00000000,
    8'b00000000,8'b00001100,8'b00011110,8'b00110011,8'b00110011,8'b00110011,8'b00000000,8'b00000000,
    8'b00000000,8'b01101110,8'b00110011,8'b00110011,8'b00110011,8'b00110011,8'b00000000,8'b00000000,
    8'b00000000,8'b00011000,8'b00101100,8'b00001100,8'b00001100,8'b00111110,8'b00001100,8'b00001000,
    8'b00000000,8'b00011111,8'b00110000,8'b00011110,8'b00000011,8'b00111110,8'b00000000,8'b00000000,
    8'b00000000,8'b00001111,8'b00000110,8'b01100110,8'b01101110,8'b00111011,8'b00000000,8'b00000000,
    8'b01111000,8'b00110000,8'b00111110,8'b00110011,8'b00110011,8'b01101110,8'b00000000,8'b00000000,
    8'b00001111,8'b00000110,8'b00111110,8'b01100110,8'b01100110,8'b00111011,8'b00000000,8'b00000000,
    8'b00000000,8'b00011110,8'b00110011,8'b00110011,8'b00110011,8'b00011110,8'b00000000,8'b00000000,
    8'b00000000,8'b00110011,8'b00110011,8'b00110011,8'b00110011,8'b00011111,8'b00000000,8'b00000000,
    8'b00000000,8'b01100011,8'b01101011,8'b01111111,8'b01111111,8'b00110011,8'b00000000,8'b00000000,
    8'b00000000,8'b00011110,8'b00001100,8'b00001100,8'b00001100,8'b00001100,8'b00001100,8'b00001110,
    8'b00000000,8'b01100111,8'b00110110,8'b00011110,8'b00110110,8'b01100110,8'b00000110,8'b00000111,
    8'b00011110,8'b00110011,8'b00110011,8'b00110000,8'b00110000,8'b00110000,8'b00000000,8'b00110000,
    8'b00000000,8'b00011110,8'b00001100,8'b00001100,8'b00001100,8'b00001110,8'b00000000,8'b00001100,
    8'b00000000,8'b01100111,8'b01100110,8'b01100110,8'b01101110,8'b00110110,8'b00000110,8'b00000111,
    8'b00011111,8'b00110000,8'b00111110,8'b00110011,8'b00110011,8'b01101110,8'b00000000,8'b00000000,
    8'b00000000,8'b00001111,8'b00000110,8'b00000110,8'b00001111,8'b00000110,8'b00110110,8'b00011100,
    8'b00000000,8'b00011110,8'b00000011,8'b00111111,8'b00110011,8'b00011110,8'b00000000,8'b00000000,
    8'b00000000,8'b01101110,8'b00110011,8'b00110011,8'b00111110,8'b00110000,8'b00110000,8'b00111000,
    8'b00000000,8'b00011110,8'b00110011,8'b00000011,8'b00110011,8'b00011110,8'b00000000,8'b00000000,
    8'b00000000,8'b00111011,8'b01100110,8'b01100110,8'b00111110,8'b00000110,8'b00000110,8'b00000111,
    8'b00000000,8'b01101110,8'b00110011,8'b00111110,8'b00110000,8'b00011110,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00011000,8'b00001100,8'b00001100,
    8'b11111111,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b01100011,8'b00110110,8'b00011100,8'b00001000,
    8'b00000000,8'b00011110,8'b00011000,8'b00011000,8'b00011000,8'b00011000,8'b00011000,8'b00011110,
    8'b00000000,8'b01000000,8'b01100000,8'b00110000,8'b00011000,8'b00001100,8'b00000110,8'b00000011,
    8'b00000000,8'b00011110,8'b00000110,8'b00000110,8'b00000110,8'b00000110,8'b00000110,8'b00011110,
    8'b00000000,8'b01111111,8'b01100110,8'b01001100,8'b00011000,8'b00110001,8'b01100011,8'b01111111,
    8'b00000000,8'b00011110,8'b00001100,8'b00001100,8'b00011110,8'b00110011,8'b00110011,8'b00110011,
    8'b00000000,8'b01100011,8'b00110110,8'b00011100,8'b00011100,8'b00110110,8'b01100011,8'b01100011,
    8'b00000000,8'b01100011,8'b01110111,8'b01111111,8'b01101011,8'b01100011,8'b01100011,8'b01100011,
    8'b00000000,8'b00001100,8'b00011110,8'b00110011,8'b00110011,8'b00110011,8'b00110011,8'b00110011,
    8'b00000000,8'b00111111,8'b00110011,8'b00110011,8'b00110011,8'b00110011,8'b00110011,8'b00110011,
    8'b00000000,8'b00011110,8'b00001100,8'b00001100,8'b00001100,8'b00001100,8'b00101101,8'b00111111,
    8'b00000000,8'b00011110,8'b00110011,8'b00111000,8'b00001110,8'b00000111,8'b00110011,8'b00011110,
    8'b00000000,8'b01100111,8'b01100110,8'b00110110,8'b00111110,8'b01100110,8'b01100110,8'b00111111,
    8'b00000000,8'b00111000,8'b00011110,8'b00111011,8'b00110011,8'b00110011,8'b00110011,8'b00011110,
    8'b00000000,8'b00001111,8'b00000110,8'b00000110,8'b00111110,8'b01100110,8'b01100110,8'b00111111,
    8'b00000000,8'b00011100,8'b00110110,8'b01100011,8'b01100011,8'b01100011,8'b00110110,8'b00011100,
    8'b00000000,8'b01100011,8'b01100011,8'b01110011,8'b01111011,8'b01101111,8'b01100111,8'b01100011,
    8'b00000000,8'b01100011,8'b01100011,8'b01101011,8'b01111111,8'b01111111,8'b01110111,8'b01100011,
    8'b00000000,8'b01111111,8'b01100110,8'b01000110,8'b00000110,8'b00000110,8'b00000110,8'b00001111,
    8'b00000000,8'b01100111,8'b01100110,8'b00110110,8'b00011110,8'b00110110,8'b01100110,8'b01100111,
    8'b00000000,8'b00011110,8'b00110011,8'b00110011,8'b00110000,8'b00110000,8'b00110000,8'b01111000,
    8'b00000000,8'b00011110,8'b00001100,8'b00001100,8'b00001100,8'b00001100,8'b00001100,8'b00011110,
    8'b00000000,8'b00110011,8'b00110011,8'b00110011,8'b00111111,8'b00110011,8'b00110011,8'b00110011,
    8'b00000000,8'b01111100,8'b01100110,8'b01110011,8'b00000011,8'b00000011,8'b01100110,8'b00111100,
    8'b00000000,8'b00001111,8'b00000110,8'b00010110,8'b00011110,8'b00010110,8'b01000110,8'b01111111,
    8'b00000000,8'b01111111,8'b01000110,8'b00010110,8'b00011110,8'b00010110,8'b01000110,8'b01111111,
    8'b00000000,8'b00011111,8'b00110110,8'b01100110,8'b01100110,8'b01100110,8'b00110110,8'b00011111,
    8'b00000000,8'b00111100,8'b01100110,8'b00000011,8'b00000011,8'b00000011,8'b01100110,8'b00111100,
    8'b00000000,8'b00111111,8'b01100110,8'b01100110,8'b00111110,8'b01100110,8'b01100110,8'b00111111,
    8'b00000000,8'b00110011,8'b00110011,8'b00111111,8'b00110011,8'b00110011,8'b00011110,8'b00001100,
    8'b00000000,8'b00011110,8'b00000011,8'b01111011,8'b01111011,8'b01111011,8'b01100011,8'b00111110,
    8'b00000000,8'b00001100,8'b00000000,8'b00001100,8'b00011000,8'b00110000,8'b00110011,8'b00011110,
    8'b00000000,8'b00000110,8'b00001100,8'b00011000,8'b00110000,8'b00011000,8'b00001100,8'b00000110,
    8'b00000000,8'b00000000,8'b00111111,8'b00000000,8'b00000000,8'b00111111,8'b00000000,8'b00000000,
    8'b00000000,8'b00011000,8'b00001100,8'b00000110,8'b00000011,8'b00000110,8'b00001100,8'b00011000,
    8'b00000110,8'b00001100,8'b00001100,8'b00000000,8'b00000000,8'b00001100,8'b00001100,8'b00000000,
    8'b00000000,8'b00001100,8'b00001100,8'b00000000,8'b00000000,8'b00001100,8'b00001100,8'b00000000,
    8'b00000000,8'b00001110,8'b00011000,8'b00110000,8'b00111110,8'b00110011,8'b00110011,8'b00011110,
    8'b00000000,8'b00011110,8'b00110011,8'b00110011,8'b00011110,8'b00110011,8'b00110011,8'b00011110,
    8'b00000000,8'b00001100,8'b00001100,8'b00001100,8'b00011000,8'b00110000,8'b00110011,8'b00111111,
    8'b00000000,8'b00011110,8'b00110011,8'b00110011,8'b00011111,8'b00000011,8'b00000110,8'b00011100,
    8'b00000000,8'b00011110,8'b00110011,8'b00110000,8'b00110000,8'b00011111,8'b00000011,8'b00111111,
    8'b00000000,8'b01111000,8'b00110000,8'b01111111,8'b00110011,8'b00110110,8'b00111100,8'b00111000,
    8'b00000000,8'b00011110,8'b00110011,8'b00110000,8'b00011100,8'b00110000,8'b00110011,8'b00011110,
    8'b00000000,8'b00111111,8'b00110011,8'b00000110,8'b00011100,8'b00110000,8'b00110011,8'b00011110,
    8'b00000000,8'b00111111,8'b00001100,8'b00001100,8'b00001100,8'b00001100,8'b00001110,8'b00001100,
    8'b00000000,8'b00111110,8'b01100111,8'b01101111,8'b01111011,8'b01110011,8'b01100011,8'b00111110,
    8'b00000000,8'b00000001,8'b00000011,8'b00000110,8'b00001100,8'b00011000,8'b00110000,8'b01100000,
    8'b00000000,8'b00001100,8'b00001100,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00111111,8'b00000000,8'b00000000,8'b00000000,
    8'b00000110,8'b00001100,8'b00001100,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00001100,8'b00001100,8'b00111111,8'b00001100,8'b00001100,8'b00000000,
    8'b00000000,8'b00000000,8'b01100110,8'b00111100,8'b11111111,8'b00111100,8'b01100110,8'b00000000,
    8'b00000000,8'b00000110,8'b00001100,8'b00011000,8'b00011000,8'b00011000,8'b00001100,8'b00000110,
    8'b00000000,8'b00011000,8'b00001100,8'b00000110,8'b00000110,8'b00000110,8'b00001100,8'b00011000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000011,8'b00000110,8'b00000110,
    8'b00000000,8'b01101110,8'b00110011,8'b00111011,8'b01101110,8'b00011100,8'b00110110,8'b00011100,
    8'b00000000,8'b01100011,8'b01100110,8'b00001100,8'b00011000,8'b00110011,8'b01100011,8'b00000000,
    8'b00000000,8'b00001100,8'b00011111,8'b00110000,8'b00011110,8'b00000011,8'b00111110,8'b00001100,
    8'b00000000,8'b00110110,8'b00110110,8'b01111111,8'b00110110,8'b01111111,8'b00110110,8'b00110110,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00110110,8'b00110110,
    8'b00000000,8'b00011000,8'b00000000,8'b00011000,8'b00011000,8'b00111100,8'b00111100,8'b00011000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,
    8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000
};

initial begin
    svp <= 0;
    hp <= 0;
    vp <= 0;
    full <= 1'b0;

    for(i = 0; i < 75; i = i + 1) begin
        for(j = 0; j < 100; j = j + 1) begin
            char_ram[i][j] <= {8{1'b0}};
        end
    end
    
    // $readmemb("font_map.txt", font_rom);
end

// TODO: offset not considered yet
assign char_vdata = vdata >> 3;
assign char_hdata = hdata >> 3;
assign valid = vdata < 600 && hdata < 800 && (full || (((char_vdata >= svp && char_vdata <= vp) ||
    ((char_vdata >= svp || char_vdata <= vp) && svp > vp)) &&
    (char_vdata != vp || char_hdata < hp)));
assign char_iv = vdata & 3'b111;
assign char_ih = hdata & 3'b111;
assign char_code = char_ram[char_vdata][char_hdata];
assign pixel = font_rom[{char_code, char_iv, char_ih}];

assign painted = valid & pixel;

assign dvi_red = {3{~painted}};
assign dvi_green = {3{~painted}};
assign dvi_blue = {2{~painted}};


reg [1:0] state;

localparam STATE_IDLE = 2'b00,
    STATE_WRITE = 2'b01;

initial begin
    state <= STATE_IDLE;
end

always @(posedge clk_bus) begin
    case(state)
        STATE_IDLE: begin
            if(cyc_i & stb_i) begin
                if(we_i) begin
                    stored_dat <= dat_i;
                    state <= STATE_WRITE;
                end
            end
        end
        STATE_WRITE: begin
            state <= STATE_IDLE;
        end
    endcase
    hp <= next_hp;
    vp <= next_vp;
    svp <= next_svp;
    full <= next_full;
    for(i = 0; i < 75; i = i + 1) begin
        for(j = 0; j < 100; j = j + 1) begin
            char_ram[i][j] <= next_char_ram[i][j];
        end
    end
end

assign ack_o = (state == STATE_WRITE);
assign next_hp = state == STATE_WRITE ? (hp == 99 ? 0 : (hp + 1)) : hp;
assign next_vp = (state == STATE_WRITE && hp == 99) ? (vp == 74 ? 0 : (vp + 1)) : vp;
assign next_svp = (state == STATE_WRITE && full) ? (svp == 74 ? 0 : (svp + 1)) : svp;
assign next_full = (state == STATE_WRITE && next_vp == svp && next_hp == 0) || 
    (state != STATE_WRITE && full);

assign rty_o = 1'b0;
assign err_o = 1'b0;

genvar ig, jg;
generate
    for(ig = 0; ig < 75; ig = ig + 1) begin
        for(jg = 0; jg < 100; jg = jg + 1) begin
            assign next_char_ram[ig][jg] = 
                state == STATE_WRITE && vp == ig && hp == jg ? stored_dat[7:0] :
                    char_ram[ig][jg];
        end
    end
endgenerate

assign de_svp = svp;
assign de_vp = vp;
assign de_hp = hp;
// assign de_valid = valid;
assign de_ascii = char_code;

endmodule